`timescale 1ns / 1ps

module Test_ALU;

	// Inputs
	reg [15:0] x;
	reg [15:0] y;
	reg zx;
	reg nx;
	reg zy;
	reg ny;
	reg f;
	reg no;

	// Outputs
	wire [15:0] out;
	wire zr;
	wire ng;

	// Instantiate the Unit Under Test (UUT)
	ALU uut (
		.x(x), 
		.y(y), 
		.zx(zx), 
		.nx(nx), 
		.zy(zy), 
		.ny(ny), 
		.f(f), 
		.no(no), 
		.out(out), 
		.zr(zr), 
		.ng(ng)
	);

	initial begin
		// Initialize Inputs
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b101010;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b111111;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b111010;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b001100;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b110000;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b001101;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b110001;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b001111;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b110011;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b011111;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b110111;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b001110;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b110010;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b010011;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b000111;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b000000;
		#100;
		x = 16'b0000000000000000;
		y = 16'b1111111111111111;
		{zx,nx,zy,ny,f,no} = 6'b010101;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b011111;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b111111;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b111010;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b001100;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b110000;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b001101;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b110001;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b001111;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b110011;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b011111;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b110111;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b001110;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b110010;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b010011;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b000111;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b000000;
		#100;
		x = 16'b0000000000010001;
		y = 16'b0000000000000011;
		{zx,nx,zy,ny,f,no} = 6'b010101;
		#100;
		// Wait 100 ns for global reset to finish
		
        
		// Add stimulus here

	end
      
endmodule

